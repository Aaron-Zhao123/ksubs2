`timescale 1ns / 1ps

//`define LOADSTORE_PORT_COUNT 0
// Kiwi Scientific Acceleration
// Start of the susbtrate for the Zynq platform.
// DRAFT !

module ksubs2_innercore(
      input 		clk,
      input 		reset_n,
      output 		led,
      output [23:0] 	pcmon,
      output reg [23:0] runtime0,
      output reg [63:0] count,
      output [23:0] 	design_serial_number,


			// Programmed I/O access to director shim
      input [7:0] 	pio_addr,
      output [31:0] 	pio_rdata,
      input [31:0] 	pio_wdata,
      input 		pio_hwen

    );
    
    wire reset;
    wire finish;
    wire [63:0] rawcount;    
    reg [1:0] controller;
    reg [23:0] runtime0_live;
    always @(posedge clk) if (!reset_n) begin
        controller <= 0;
	runtime0 <= 0;
	runtime0_live <= 0;
	count <= 101; // for debug
        end
        else begin
	     count <= rawcount;
             if (controller == 0) begin
	     	      controller <= 1;
		      runtime0_live <= 0;
		      runtime0 <= runtime0_live;
		      end
             if (controller == 1) controller <= 2;
             if (controller == 2 && runtime0_live != 24'hffffff) runtime0_live <= runtime0_live + 1; 
             if (controller == 2 && finished) controller <= 3; 
             if (controller == 3) controller <= 0;
             end
             
    assign kreset = (controller == 0);
    parameter dram_dwidth = 256;          // 32 byte DRAM burst size or cache line.
    parameter laneSize = 8;
    parameter noLanes = dram_dwidth / laneSize; // Bytelanes.
    parameter memsize = 64;
 
    wire [noLanes-1:0] bs_r0bank_lanes;
    wire [21:0]         bs_r0bank_addr;
    wire bs_r0bank_oprdy, bs_r0bank_opreq, bs_r0bank_ack, bs_r0bank_rwbar;
    wire [dram_dwidth-1:0]  bs_r0bank_rdata, bs_r0bank_wdata;
 
    wire [noLanes-1:0] fs_r0bank_lanes;
    wire [21:0]         fs_r0bank_addr;
    wire fs_r0bank_oprdy, fs_r0bank_opreq, fs_r0bank_ack, fs_r0bank_rwbar;
    wire [dram_dwidth-1:0]  fs_r0bank_rdata, fs_r0bank_wdata;
    
  

   // The design of interest - generated by KiwiC or otherwise.
    up_counter dut(.clk(clk), 
		       .reset(kreset),

// old director interface
//		.pcmon(pcmon),
		       .led(led),
		       .finished(finished),
		       .count(rawcount),
		       .design_serial_number(design_serial_number),

/*
`ifdef LOADSTORE_PORT_COUNT
		       // connect 'off-chip' memory to BRAM for now
		       .hf1_dram0bank_lanes(fs_r0bank_lanes),
		       .hf1_dram0bank_oprdy(fs_r0bank_oprdy),
		       .hf1_dram0bank_opreq(fs_r0bank_opreq),
		       .hf1_dram0bank_ack(fs_r0bank_ack),
		       .hf1_dram0bank_rwbar(fs_r0bank_rwbar),   .hf1_dram0bank_rdata(fs_r0bank_rdata),
		       .hf1_dram0bank_addr(fs_r0bank_addr),     .hf1_dram0bank_wdata(fs_r0bank_wdata),
`endif
*/
		       // Programmed I/O access to director shim
		       .pio_hwen(pio_hwen), .pio_rdata(pio_rdata), .pio_wdata(pio_wdata), .pio_addr(pio_addr)
		       
    );

/*
`ifdef LOADSTORE_PORT_COUNT
   membank256_hf1    #(noLanes, laneSize, memsize) drambank0_hfast1
   		  (clk, reset,
		      fs_r0bank_rwbar, fs_r0bank_rdata,
		      fs_r0bank_wdata, fs_r0bank_addr,
		      fs_r0bank_oprdy, fs_r0bank_opreq,
		      fs_r0bank_ack, fs_r0bank_lanes);
`endif
  */ 
endmodule
